library verilog;
use verilog.vl_types.all;
entity Lab3_Part1_vlg_vec_tst is
end Lab3_Part1_vlg_vec_tst;
